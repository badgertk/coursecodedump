** Part 1 - Current Mirror - AC Analysis **
.INCLUDE sedra_lib.lib

* DC and AC Sources
VD VDD 0 DC 3.3V AC 1
V1 D1 0 DC 1.0883V
V2 D2 0 DC 1.0883V

* Resistors
R VDD D0 23.541K

* MOSFETs
M0 D0 D0 0 0 NMOS0P5 W=5U L=0.5U
M1 D1 D0 0 0 NMOS0P5 W=50U L=0.5U
M2 D2 D0 0 0 NMOS0P5 W=250U L=0.5U

** AC Analysis
.OPTIONS POST
.OP
.AC DEC 10 1 1E6

.END
